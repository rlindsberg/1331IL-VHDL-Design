-- WIP
library ieee;
use ieee.std_logic_1164.all;

entity b8_carry_select_adder is
	port(
		);
end entity;

architecture gooy_inside of b8_carry_select_adder is
	component full_adder
end architecture;