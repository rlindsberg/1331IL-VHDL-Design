Entity enchip is
  Port( clk     :     std_logic;
        reset   :     std_logic;
        stop    :     std_logic;
        choice  :     std_logic;
        s       : out std_logic_vector(3 downto 0));
End Entity;

Architecture structure of enchip is
  
End Architecture;
