entity adder is
  port (
    a   : std_logica_vector(7 downto 0);
    b   : std_logica_vector(7 downto 0);
    sum : out std_logica_vector(7 downto 0)
  );
end entity;
