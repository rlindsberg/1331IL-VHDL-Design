Entity ROM is
  Port(
    addr: in address_bus;
    data: out instruction_bus;
    ce: in std_logic
  );
End;

Architecture behavioural of ROM is
  Signal
  Begin
    Process
      Begin

End behavioural;
