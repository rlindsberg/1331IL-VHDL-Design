entity Adder is
  port(
    a : unsigned(7 downto 0);
    b : unsigned(7 downto 0)

  )
