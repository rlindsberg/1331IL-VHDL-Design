Entity DataBuffer is
  Port(
    out_en: in std_logic;
    data_in: in data_word;
    data_out: out data_bus
  );
End;

Architecture behavioural of DataBuffer is

  Signal

Begin

End behavioural;
